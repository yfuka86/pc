0:10,346,3.46
1:10,392,3.92
2:15,615,2.73333
3:16,846,3.30469
4:19,1696,4.69806
5:20,1159,2.8975
6:20,1443,3.6075
7:20,1393,3.4825
8:20,1377,3.4425
9:25,2458,3.9328
10:27,2168,2.97394
11:30,2679,2.97667
12:30,2550,2.83333
13:30,2436,2.70667
14:35,3927,3.20571
15:40,4015,2.50937
16:40,3241,2.02562
17:50,6316,2.5264
18:50,4359,1.7436
19:100,11027,1.1027
0:10,360,3.6
1:10,345,3.45
2:15,775,3.44444
3:16,1268,4.95312
4:19,1599,4.42936
5:20,1388,3.47
6:20,1665,4.1625
7:20,1775,4.4375
8:20,1359,3.3975
9:25,2701,4.3216
10:27,2000,2.74348
11:30,2339,2.59889
12:30,2099,2.33222
13:30,2494,2.77111
14:35,3934,3.21143
15:40,4057,2.53563
16:40,3289,2.05563
17:50,6489,2.5956
18:50,4334,1.7336
19:100,10984,1.0984
0:10,289,2.89
1:10,464,4.64
2:15,786,3.49333
3:16,855,3.33984
4:19,1680,4.65374
5:20,1531,3.8275
6:20,1734,4.335
7:20,1499,3.7475
8:20,1489,3.7225
9:25,2438,3.9008
10:27,2265,3.107
11:30,2517,2.79667
12:30,2224,2.47111
13:30,2405,2.67222
14:35,3838,3.13306
15:40,4024,2.515
16:40,3209,2.00563
17:50,6436,2.5744
18:50,4364,1.7456
19:100,11045,1.1045
0:10,300,3
1:10,430,4.3
2:15,762,3.38667
3:16,814,3.17969
4:19,1494,4.1385
5:20,1201,3.0025
6:20,1511,3.7775
7:20,1443,3.6075
8:20,1392,3.48
9:25,2656,4.2496
10:27,2325,3.1893
11:30,2708,3.00889
12:30,2276,2.52889
13:30,2541,2.82333
14:35,3730,3.0449
15:40,4087,2.55437
16:40,3256,2.035
17:50,6397,2.5588
18:50,4358,1.7432
19:100,11029,1.1029
0:10,304,3.04
1:10,347,3.47
2:15,804,3.57333
3:16,855,3.33984
4:19,1596,4.42105
5:20,1158,2.895
6:20,1488,3.72
7:20,1827,4.5675
8:20,1432,3.58
9:25,2343,3.7488
10:27,2220,3.04527
11:30,2578,2.86444
12:30,2102,2.33556
13:30,2468,2.74222
14:35,3758,3.06776
15:40,4043,2.52687
16:40,3195,1.99687
17:50,6386,2.5544
18:50,4439,1.7756
19:100,10968,1.0968
